// Code your testbench here
// or browse Examples
`include "testbench_top.sv"     